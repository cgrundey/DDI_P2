////////////////////////////////////////////////////////////////////////////////
// Filename:    tb_register12bit_cgrundey.v
// Author:      Colin Grundey
// Date:        19 March 2018
// Version:     1
// Description: Test bench for 12-bit register implementation
////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/100ps

module tb_register12bit_cgrundey();

	initial begin

	end

endmodule
